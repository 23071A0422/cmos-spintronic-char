magic
tech sky130A
timestamp 1704283200
<< nwell >>
rect 0 80 100 160
<< pdiffusion >>
rect 10 90 90 150
<< ndiffusion >>
rect 10 10 90 70
<< polysilicon >>
rect 45 5 55 155
<< metal1 >>
rect 0 150 100 160 ;# VDD Rail
rect 0 0 100 10 ;# GND Rail
rect 40 75 60 85 ;# Output Pin
<< labels >>
label vdd 50 155
label gnd 50 5
label in 50 10
label out 50 80